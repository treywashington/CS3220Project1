module SetClock(OUT,IN);

endmodule